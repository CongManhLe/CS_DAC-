* Extracted by KLayout with SG13G2 LVS runset on : 22/01/2026 23:57

.SUBCKT inverter VSS VDD Y A
M$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 VDD A Y VDD sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS inverter
