** sch_path: /home/lecongmanh/CS_DAC/xschem/Test_thermo.sch
**.subckt Test_thermo
x3 D1 D2 D3 D4 D5 D6 D7 X5 X6 X7 VDD VSS thermo_decoder
V8 X5 GND PULSE(0 1 0 5n 5n 795n 1600n)
V9 X6 GND PULSE(0 1 0 5n 5n 1595n 3200n)
V13 X7 GND PULSE(0 1 0 5n 5n 3195n 6400n)
V1 VDD GND 1
V2 VSS GND 0
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerDIO.lib dio_tt
.include /home/lecongmanh/unic-cass/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice





.save v(D1) v(D2) v(D3) v(D4) v(D5) v(D6) v(D7)
.control
.options method=gear
set wr_vecnames
set wr_singlescale
tran 0.1n 6400n
run
plot v(D1) v(D2) v(D3) v(D4) v(D5) v(D6) v(D7)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  thermo_decoder.sym # of pins=12
** sym_path: /home/lecongmanh/CS_DAC/xschem/thermo_decoder.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/thermo_decoder.sch
.subckt thermo_decoder D1 D2 D3 D4 D5 D6 D7 X0 X1 X2 VDD VSS
*.ipin X2
*.ipin X1
*.ipin X0
*.opin D7
*.opin D6
*.opin D5
*.opin D4
*.opin D3
*.opin D1
*.opin D2
*.ipin VDD
*.ipin VSS
x1 net1 X1 X0 VDD VSS sg13g2_and2_2
x2 D7 X2 net1 VDD VSS sg13g2_and2_2
x3 D6 X1 X2 VDD VSS sg13g2_and2_2
x4 D2 X2 X1 VDD VSS sg13g2_or2_2
x5 D1 X0 D2 VDD VSS sg13g2_or2_2
x6 net2 X0 X1 VDD VSS sg13g2_or2_2
x7 D5 net2 X2 VDD VSS sg13g2_and2_2
x8 net3 X0 X1 VDD VSS sg13g2_and2_2
x9 D3 net3 X2 VDD VSS sg13g2_or2_2
x10 D4 X2 VDD VSS sg13g2_buf_2
.ends

.GLOBAL GND
.end
