** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_DAC_10b_test.sch
**.subckt CS_DAC_10b_test
V1 VDD GND 1
V3 VBIAS GND 1
V2 CLK GND PULSE(0 1 0n 5n 5n 20n 50n)
V4 X1 GND PULSE(0 1 0 5n 5n 45n 100n)
V5 X2 GND PULSE(0 1 0 5n 5n 95n 200n)
V6 X3 GND PULSE(0 1 0 5n 5n 195n 400n)
V7 X4 GND PULSE(0 1 0 5n 5n 395n 800n)
V8 X5 GND PULSE(0 1 0 5n 5n 795n 1600n)
V9 X6 GND PULSE(0 1 0 5n 5n 1595n 3200n)
x4 CLK OUTN OUTP VBIAS VDD GND X1 X10 X2 X3 X4 X5 X6 X7 X8 X9 CS_DAC_10b
V13 X7 GND PULSE(0 1 0 5n 5n 3195n 6400n)
V15 X8 GND PULSE(0 1 0 5n 5n 6395n 12800n)
V17 X9 GND PULSE(0 1 0 1n 1n 12795n 25600n)
V19 X10 GND PULSE(0 1 0 1n 1n 25595n 51200n)
Vds net1 GND 1.5
Vd net1 OUTN 0
.save i(vd)
Vd1 net1 OUTP 0
.save i(vd1)
**** begin user architecture code


.save i(Vd) i(Vd1)
.control
.options method=gear
set wr_vecnames
set wr_singlescale
tran 0.1n 51200n
run
write CS_DAC_10b.raw i(Vd) i(Vd1)
.endc





.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerDIO.lib dio_tt
.include /home/lecongmanh/unic-cass/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



**** end user architecture code
**.ends

* expanding   symbol:  CS_DAC_10b.sym # of pins=16
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_DAC_10b.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_DAC_10b.sch
.subckt CS_DAC_10b CLK OUTN OUTP VBIAS VDD VSS X1 X10 X2 X3 X4 X5 X6 X7 X8 X9
*.ipin X9
*.ipin X8
*.ipin X7
*.ipin X6
*.ipin X5
*.ipin X4
*.ipin X3
*.ipin X2
*.ipin X10
*.ipin X1
*.iopin VSS
*.ipin VDD
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin CLK
x1 net8 net9 net10 net11 net12 net13 net14 CLK net1 net2 net3 net4 net5 net6 net7 OUTN OUTP VBIAS VDD VSS 6MSB
x2 CLK OUTN OUTP VBIAS VDD VSS X1 X2 X3 X4 4MSB_weighted
x3 net8 net9 net10 net11 net12 net13 net14 X5 X6 X7 VDD VSS thermo_decoder
x5 net1 net2 net3 net4 net5 net6 net7 X8 X9 X10 VDD VSS thermo_decoder
.ends


* expanding   symbol:  6MSB.sym # of pins=20
** sym_path: /home/lecongmanh/CS_DAC/xschem/6MSB.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/6MSB.sch
.subckt 6MSB C1 C2 C3 C4 C5 C6 C7 CLK D1 D2 D3 D4 D5 D6 D7 OUTN OUTP VBIAS VDD VSS
*.iopin VSS
*.ipin VDD
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin D7
*.ipin D6
*.ipin D5
*.ipin D4
*.ipin D3
*.ipin D2
*.ipin D1
*.ipin CLK
*.ipin C7
*.ipin C6
*.ipin C5
*.ipin C4
*.ipin C3
*.ipin C2
*.ipin C1
x33 CLK C1 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x1 CLK C2 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x2 CLK C3 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x3 CLK C4 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x4 CLK C5 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x5 CLK C6 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x6 CLK C7 OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x7 CLK VSS OUTN OUTP D1 VDD VBIAS VDD VSS Unit_cell
x8 CLK C1 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x9 CLK C2 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x10 CLK C3 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x11 CLK C4 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x12 CLK C5 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x13 CLK C6 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x14 CLK C7 OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x15 CLK VSS OUTN OUTP D2 D1 VBIAS VDD VSS Unit_cell
x16 CLK C1 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x17 CLK C2 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x18 CLK C3 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x19 CLK C4 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x20 CLK C5 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x21 CLK C6 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x22 CLK C7 OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x23 CLK VSS OUTN OUTP D3 D2 VBIAS VDD VSS Unit_cell
x24 CLK C1 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x25 CLK C2 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x26 CLK C3 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x27 CLK C4 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x28 CLK C5 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x29 CLK C6 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x30 CLK C7 OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x31 CLK VSS OUTN OUTP D4 D3 VBIAS VDD VSS Unit_cell
x32 CLK C1 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x34 CLK C2 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x35 CLK C3 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x36 CLK C4 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x37 CLK C5 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x38 CLK C6 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x39 CLK C7 OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x40 CLK VSS OUTN OUTP D5 D4 VBIAS VDD VSS Unit_cell
x41 CLK C1 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x42 CLK C2 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x43 CLK C3 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x44 CLK C4 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x45 CLK C5 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x46 CLK C6 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x47 CLK C7 OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x48 CLK VSS OUTN OUTP D6 D5 VBIAS VDD VSS Unit_cell
x49 CLK C1 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x50 CLK C2 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x51 CLK C3 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x52 CLK C4 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x53 CLK C5 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x54 CLK C6 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x55 CLK C7 OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x56 CLK VSS OUTN OUTP D7 D6 VBIAS VDD VSS Unit_cell
x57 CLK C1 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x58 CLK C2 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x59 CLK C3 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x60 CLK C4 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x61 CLK C5 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x62 CLK C6 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
x63 CLK C7 OUTN OUTP VSS D7 VBIAS VDD VSS Unit_cell
.ends


* expanding   symbol:  4MSB_weighted.sym # of pins=10
** sym_path: /home/lecongmanh/CS_DAC/xschem/4MSB_weighted.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/4MSB_weighted.sch
.subckt 4MSB_weighted CLK OUTN OUTP VBIAS VDD VSS X1 X2 X3 X4
*.ipin X4
*.ipin X3
*.ipin X2
*.ipin X1
*.iopin VSS
*.ipin VDD
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin CLK
x9 net2 net1 OUTN OUTP VBIAS VSS CS_Switch_1x
x2 net4 net3 OUTN OUTP VBIAS VSS CS_Switch_2x
x3 net6 net5 OUTN OUTP VBIAS VSS CS_Switch_4x
x5 net8 net7 OUTN OUTP VBIAS VSS CS_Switch_8x
x1 net1 net2 CLK X1 VDD VDD VSS sg13g2_dfrbp_2
x4 net3 net4 CLK X2 VDD VDD VSS sg13g2_dfrbp_2
x6 net5 net6 CLK X3 VDD VDD VSS sg13g2_dfrbp_2
x7 net7 net8 CLK X4 VDD VDD VSS sg13g2_dfrbp_2
.ends


* expanding   symbol:  thermo_decoder.sym # of pins=12
** sym_path: /home/lecongmanh/CS_DAC/xschem/thermo_decoder.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/thermo_decoder.sch
.subckt thermo_decoder D1 D2 D3 D4 D5 D6 D7 X0 X1 X2 VDD VSS
*.ipin X2
*.ipin X1
*.ipin X0
*.opin D7
*.opin D6
*.opin D5
*.opin D4
*.opin D3
*.opin D1
*.opin D2
*.ipin VDD
*.ipin VSS
x1 net1 X1 X0 VDD VSS sg13g2_and2_2
x2 D7 X2 net1 VDD VSS sg13g2_and2_2
x3 D6 X1 X2 VDD VSS sg13g2_and2_2
x4 D2 X2 X1 VDD VSS sg13g2_or2_2
x5 D1 X0 D2 VDD VSS sg13g2_or2_2
x6 net2 X0 X1 VDD VSS sg13g2_or2_2
x7 D5 net2 X2 VDD VSS sg13g2_and2_2
x8 net3 X0 X1 VDD VSS sg13g2_and2_2
x9 D3 net3 X2 VDD VSS sg13g2_or2_2
x10 D4 X2 VDD VSS sg13g2_buf_2
.ends


* expanding   symbol:  Unit_cell.sym # of pins=9
** sym_path: /home/lecongmanh/CS_DAC/xschem/Unit_cell.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/Unit_cell.sch
.subckt Unit_cell CLK Ci OUTN OUTP Ri Ri-1 VBIAS VDD VSS
*.iopin VSS
*.ipin VDD
*.ipin VBIAS
*.ipin Ri-1
*.ipin Ri
*.iopin OUTP
*.iopin OUTN
*.ipin Ci
*.ipin CLK
x1 net5 net4 OUTN OUTP VBIAS VSS CS_Switch_16x
x2 net1 Ri Ci VDD VSS sg13g2_or2_2
x3 net6 net1 Ri-1 VDD VSS sg13g2_nand2_2
x6 net2 net3 CLK net7 VDD VDD VSS sg13g2_dfrbp_2
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
x4 net4 net2 VDD VSS sg13g2_buf_2
x5 net5 net3 VDD VSS sg13g2_buf_2
x7 net7 net6 VDD VSS sg13g2_buf_2
.ends


* expanding   symbol:  CS_Switch_1x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_1x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_1x.sch
.subckt CS_Switch_1x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM6 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM1 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM8 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM9 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM10 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM11 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM12 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM3 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM4 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM13 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM14 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM15 VSS VSS VSS VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
.ends


* expanding   symbol:  CS_Switch_2x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_2x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_2x.sch
.subckt CS_Switch_2x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=0.6u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=0.6u l=0.45u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends


* expanding   symbol:  CS_Switch_4x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_4x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_4x.sch
.subckt CS_Switch_4x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=1.2u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=1.2u l=0.45u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends


* expanding   symbol:  CS_Switch_8x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_8x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_8x.sch
.subckt CS_Switch_8x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=2.4u l=0.48u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=2.4u l=0.48u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends


* expanding   symbol:  CS_Switch_16x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_16x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_16x.sch
.subckt CS_Switch_16x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=5.2u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=5.2u l=0.45u ng=1 m=1
C2 net1 GND 1u m=1
.ends

.GLOBAL GND
.end
