* Extracted by KLayout with SG13G2 LVS runset on : 22/01/2026 22:49

.SUBCKT TOP
M$1 \$3 A Y \$1 sg13_lv_nmos L=0.135u W=0.15u AS=0.1005p AD=0.09975p PS=1.34u
+ PD=1.33u
M$2 VDD A Y VDD sg13_lv_pmos L=0.135u W=0.15u AS=0.1005p AD=0.09975p PS=1.34u
+ PD=1.33u
.ENDS TOP
