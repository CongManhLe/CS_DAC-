** sch_path: /home/lecongmanh/CS_DAC/xschem/4LSB_Test.sch
**.subckt 4LSB_Test
x2 CLK net1 net2 VBIAS VDD VSS X1 X2 X3 X4 4MSB_weighted
V1 VDD GND 1
V3 VBIAS GND 1
V2 CLK GND PULSE(0 1 0n 5n 5n 20n 50n)
V4 X1 GND PULSE(0 1 0 5n 5n 45n 100n)
V5 X2 GND PULSE(0 1 0 5n 5n 95n 200n)
V6 X3 GND PULSE(0 1 0 5n 5n 195n 400n)
V7 X4 GND PULSE(0 1 0 5n 5n 395n 800n)
V8 VSS GND 0
Vds net3 GND 1.5
Vd net3 net1 0
.save i(vd)
Vd1 net3 net2 0
.save i(vd1)
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ
.lib cornerDIO.lib dio_tt
.include /home/lecongmanh/unic-cass/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice





.save i(Vd) i(Vd1)
.control
.options method=gear
set wr_vecnames
set wr_singlescale
tran 0.1n 1600n
run
write 4LSB.raw i(Vd) i(Vd1)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  4MSB_weighted.sym # of pins=10
** sym_path: /home/lecongmanh/CS_DAC/xschem/4MSB_weighted.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/4MSB_weighted.sch
.subckt 4MSB_weighted CLK OUTN OUTP VBIAS VDD VSS X1 X2 X3 X4
*.ipin X4
*.ipin X3
*.ipin X2
*.ipin X1
*.iopin VSS
*.ipin VDD
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin CLK
x9 net2 net1 OUTN OUTP VBIAS VSS CS_Switch_1x
x2 net4 net3 OUTN OUTP VBIAS VSS CS_Switch_2x
x3 net6 net5 OUTN OUTP VBIAS VSS CS_Switch_4x
x5 net8 net7 OUTN OUTP VBIAS VSS CS_Switch_8x
x1 net1 net2 CLK X1 VDD VDD VSS sg13g2_dfrbp_2
x4 net3 net4 CLK X2 VDD VDD VSS sg13g2_dfrbp_2
x6 net5 net6 CLK X3 VDD VDD VSS sg13g2_dfrbp_2
x7 net7 net8 CLK X4 VDD VDD VSS sg13g2_dfrbp_2
.ends


* expanding   symbol:  CS_Switch_1x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_1x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_1x.sch
.subckt CS_Switch_1x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM6 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM1 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM8 OUTP INP net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM9 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM10 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM11 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM12 OUTN INN net1 VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM3 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM4 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM13 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM14 net1 VSS VSS VSS sg13_lv_nmos w=0.5u l=0.13u ng=1 m=1
XM15 VSS VSS VSS VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
.ends


* expanding   symbol:  CS_Switch_2x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_2x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_2x.sch
.subckt CS_Switch_2x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=0.6u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=0.6u l=0.45u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends


* expanding   symbol:  CS_Switch_4x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_4x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_4x.sch
.subckt CS_Switch_4x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=1.2u l=0.45u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=1.2u l=0.45u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends


* expanding   symbol:  CS_Switch_8x.sym # of pins=6
** sym_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_8x.sym
** sch_path: /home/lecongmanh/CS_DAC/xschem/CS_Switch_8x.sch
.subckt CS_Switch_8x INN INP OUTN OUTP VBIAS VSS
*.iopin VSS
*.ipin VBIAS
*.iopin OUTP
*.iopin OUTN
*.ipin INP
*.ipin INN
XM1 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 OUTP INP net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM3 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM4 OUTN INN net1 VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM7 net1 VBIAS net2 VSS sg13_hv_nmos w=2.4u l=0.48u ng=1 m=1
XM5 net2 VBIAS VSS VSS sg13_hv_nmos w=2.4u l=0.48u ng=1 m=1
C1 OUTP GND 1u m=1
C2 OUTN GND 1u m=1
C3 net1 GND 1u m=1
.ends

.GLOBAL GND
.end
